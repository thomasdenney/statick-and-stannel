`include "defaults.vh"

`define CORE_MESSAGE_NONE            4'd15
`define CORE_MESSAGE_START_PROCESS   `OP_PROCESS_START
`define CORE_MESSAGE_YIELD           `OP_PROCESS_YIELD
`define CORE_MESSAGE_HALT            `OP_PROCESS_END
`define CORE_MESSAGE_CREATE_CHANNEL  `OP_PROCESS_CREATE_CHANNEL
`define CORE_MESSAGE_DELETE_CHANNEL  `OP_PROCESS_DESTROY_CHANNEL
`define CORE_MESSAGE_SEND            `OP_PROCESS_SEND
`define CORE_MESSAGE_RECEIVE         `OP_PROCESS_RECEIVE
`define CORE_MESSAGE_ALT_START       `OP_PROCESS_ALT_START
`define CORE_MESSAGE_ALT_WAIT        `OP_PROCESS_ALT_WAIT
`define CORE_MESSAGE_ALT_END         `OP_PROCESS_ALT_END
`define CORE_MESSAGE_ENABLE_CHANNEL  `OP_PROCESS_ENABLE_CHANNEL
`define CORE_MESSAGE_DISABLE_CHANNEL `OP_PROCESS_DISABLE_CHANNEL

`define PROCESSOR_MESSAGE_NONE                        3'd0
`define PROCESSOR_MESSAGE_RESUME                      3'd1
`define PROCESSOR_MESSAGE_RECEIVE                     3'd2
`define PROCESSOR_MESSAGE_RECEIVE_AND_JUMP            3'd3
`define PROCESSOR_MESSAGE_RECEIVE_AND_JUMP_AND_WAIT   3'd4
`define PROCESSOR_MESSAGE_RESUME_AND_WAIT             3'd5
