// Baud rates. These are derived from dividing 12,000,000 Hz by the
// target rate and then rounding down.
`define B115200 104