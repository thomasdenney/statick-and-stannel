`define REG_PC  3'b000
`define REG_SP  3'b001
`define REG_CSP 3'b010
`define REG_S1  3'b011
`define REG_S2  3'b100
`define REG_S3  3'b101